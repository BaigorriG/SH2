library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.HexaPackage.all;

ENTITY CONTROLADOR_VGA IS
	GENERIC( BITS:	INTEGER:=10);
	PORT(
		CLK			:	IN	STD_LOGIC;
		CLR			:	IN	STD_LOGIC;
		RED_IN		:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		GREEN_IN		:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLUE_IN		:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		
		HSYNC			:	OUT	STD_LOGIC;
		VSYNC			:	OUT	STD_LOGIC;
		VGA_SYNC_N	:	OUT	STD_LOGIC;
		VGA_BLANK_N	:	OUT	STD_LOGIC;
		X				:	OUT	UNSIGNED(BITS-1 DOWNTO 0);
		Y				:	OUT	UNSIGNED(BITS-1 DOWNTO 0);
		RED			:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		GREEN			:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLUE			:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		END_FRAME	:	OUT	STD_LOGIC;
		PRE_FRAME	:	OUT	STD_LOGIC
		);
END ENTITY;

ARCHITECTURE BEH OF CONTROLADOR_VGA IS


CONSTANT HPIXELS	: UNSIGNED:= TO_UNSIGNED(800,BITS);		--SYNC_PULSE	+BP	+AREA VISIBLE	+FP
CONSTANT vLINES	: UNSIGNED:= TO_UNSIGNED(525,BITS);
CONSTANT HPULSE	: UNSIGNED:= TO_UNSIGNED(96,BITS);				--96
CONSTANT VPULSE	: UNSIGNED:= TO_UNSIGNED(2,BITS);				--2
CONSTANT HBP		: UNSIGNED:= TO_UNSIGNED(144,BITS);							--48
CONSTANT VBP		: UNSIGNED:= TO_UNSIGNED(35,BITS);								--33
CONSTANT HAREA		: UNSIGNED:= TO_UNSIGNED(640,BITS);									--640
CONSTANT VAREA		: UNSIGNED:= TO_UNSIGNED(480,BITS);									--480
CONSTANT HFP		: UNSIGNED:= TO_UNSIGNED(784,BITS);														--16
CONSTANT VFP		: UNSIGNED:= TO_UNSIGNED(515,BITS);														--10

----PARA PROBAR 800X600 -- SE NECESITA GENERAR RELOJ DE 40 MHZ
--
--CONSTANT HPIXELS	: UNSIGNED:= TO_UNSIGNED(1056,BITS);		--SYNC_PULSE	+BP	+AREA VISIBLE	+FP
--CONSTANT vLINES	: UNSIGNED:= TO_UNSIGNED(628,BITS);
--CONSTANT HPULSE	: UNSIGNED:= TO_UNSIGNED(128,BITS);				--128
--CONSTANT VPULSE	: UNSIGNED:= TO_UNSIGNED(4,BITS);					--4
--CONSTANT HBP		: UNSIGNED:= TO_UNSIGNED(216,BITS);						--88
--CONSTANT VBP		: UNSIGNED:= TO_UNSIGNED(27,BITS);						--23
--CONSTANT HAREA		: UNSIGNED:= TO_UNSIGNED(800,BITS);									--800
--CONSTANT VAREA		: UNSIGNED:= TO_UNSIGNED(600,BITS);									--600
--CONSTANT HFP		: UNSIGNED:= TO_UNSIGNED(1016,BITS);													--40
--CONSTANT VFP		: UNSIGNED:= TO_UNSIGNED(627,BITS);													--1



SIGNAL	HC	:	UNSIGNED(BITS-1 DOWNTO 0);
SIGNAL	VC	:	UNSIGNED(BITS-1 DOWNTO 0);
SIGNAL	IN_FRAME	:	STD_LOGIC;
SIGNAL 	VGA_SYNC,VGA_BLANK:	STD_LOGIC;
BEGIN

HSYNC<='0' WHEN (HC<HPULSE) ELSE '1';
VSYNC<='0' WHEN (VC<VPULSE) ELSE '1';
VGA_SYNC	<= '1' WHEN	(VC >= VBP AND VC < VFP) ELSE '0';
VGA_BLANK<=	'1' WHEN (HC >= HBP AND HC < HFP) ELSE '0';
IN_FRAME <= '1' WHEN (VGA_SYNC='1' AND VGA_BLANK='1') ELSE '0';
PRE_FRAME <= '1' WHEN (HC=(BITS-1 DOWNTO 0 => '0') AND VC=(BITS-1 DOWNTO 0 => '0')) ELSE '0';
END_FRAME <= '1' WHEN (HC=(BITS-1 DOWNTO 0 => '0') AND VC=VFP) ELSE '0';

VGA_BLANK_N<=VGA_BLANK;
VGA_SYNC_N<=VGA_SYNC;

SUMACONTADORES:PROCESS (CLK,CLR,HC,VC)
BEGIN
IF (CLR='1') THEN
	HC<=(OTHERS=>'0');
	VC<=(OTHERS=>'0');
ELSIF (RISING_EDGE(CLK)) THEN

	IF(HC < HPIXELS-1) THEN
		HC<=HC+1;
	ELSE
		HC<=(OTHERS=>'0');
		IF(VC < VLINES-1) THEN
			VC<=VC+1;
		ELSE
			VC<=(OTHERS=>'0');
		END IF;
	END IF;
END IF;
END PROCESS;

SETEACOORDENADAS:PROCESS (CLK)
BEGIN
	IF(RISING_EDGE(CLK)) THEN
		IF(VC >= VBP AND VC < VFP) THEN
			Y <= VC-VBP;
		ELSE
			Y <= (OTHERS=>'0');
		END IF;
		IF(HC >= HBP AND HC < HFP) THEN
			X <= HC-HBP;
		ELSE
			X	<=	(OTHERS=>'0');
		END IF;
	END IF;
END PROCESS;

SETEACOLORES:PROCESS (CLK)
BEGIN
IF RISING_EDGE(CLK) THEN
	IF (IN_FRAME='1') THEN
		RED <= RED_IN;
		GREEN <= GREEN_IN;
		BLUE <= BLUE_IN;
	ELSE
		RED <= (OTHERS => '0');
		GREEN <= (OTHERS => '0');
		BLUE <= (OTHERS => '0');
	END IF;
END IF;
END PROCESS;

END ARCHITECTURE;
