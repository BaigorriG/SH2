library ieee; 
use ieee.std_logic_1164.all;

ENTITY DATA_BUFFER IS
GENERIC(
			data_width:	integer:=8
		);
PORT(
	DATAIN:	IN		STD_LOGIC_VECTOR(data_width-1 DOWNTO 0);
	EN:		IN		STD_LOGIC;
	CLK:		IN		STD_LOGIC;
	CLEAR:	IN		STD_LOGIC;
	DATAOUT:	OUT	STD_LOGIC_VECTOR(data_width-1 DOWNTO 0)
	);
END DATA_BUFFER;

ARCHITECTURE BEH OF DATA_BUFFER IS

BEGIN
STORE: PROCESS	(CLK,EN,CLEAR)
BEGIN
	IF (CLEAR='1') THEN
		DATAOUT<=(OTHERS=>'0');
	ELSIF (RISING_EDGE(CLK) AND EN='1') THEN
		DATAOUT<=DATAIN;
	END IF;
END PROCESS;
END BEH;