library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE HexaPackage IS

CONSTANT BITS		: INTEGER:=	10;
function bit2bool(b: std_logic) return boolean;
CONSTANT CENTROX	: SIGNED:= TO_SIGNED(320,BITS);
CONSTANT CENTROY	: SIGNED:= TO_SIGNED(240,BITS);

--------------------------------------------------------------------------------------------------------------------
----------------------------------------------COMPONENTES-----------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------

COMPONENT PLL IS
	PORT
	(
		areset		: IN STD_LOGIC  := '0';
		inclk0		: IN STD_LOGIC  := '0';
		c0		: OUT STD_LOGIC 
	);
END COMPONENT;

COMPONENT CONTROLADOR_VGA IS
	GENERIC( BITS:	INTEGER:=10);
	PORT(
		CLK			:	IN	STD_LOGIC;
		CLR			:	IN	STD_LOGIC;
		RED_IN		:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		GREEN_IN		:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLUE_IN		:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		
		HSYNC			:	OUT	STD_LOGIC;
		VSYNC			:	OUT	STD_LOGIC;
		VGA_SYNC_N	:	OUT	STD_LOGIC;
		VGA_BLANK_N	:	OUT	STD_LOGIC;
		X				:	OUT	UNSIGNED(BITS-1 DOWNTO 0);
		Y				:	OUT	UNSIGNED(BITS-1 DOWNTO 0);
		RED			:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		GREEN			:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLUE			:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		END_FRAME	:	OUT	STD_LOGIC;
		PRE_FRAME	:	OUT	STD_LOGIC
		);
END COMPONENT;

component DesplazaXYalCentro is

	port(
		Clk		:	in	std_logic;
		Xin		:	in unsigned(9 downto 0);
		Yin		:	in unsigned(9 downto 0);
		Xout		:	out signed(9 downto 0);
		Yout		:	out signed(9 downto 0)
	);
end component;

component rotar is
	port(
		clk			:	in std_logic;
		Actualizar	:	in std_logic;
		X_in			:	in signed(9 downto 0);
		Y_in			:	in signed(9 downto 0);
		angulo		:	in	unsigned(9 downto 0);
		
		X_out			:	out	signed(9 downto 0);
		Y_out			:	out	signed(9 downto 0)
	);
end component;

component conv_hexagonal is
	port(
		clk			: in std_logic;
		x				: in signed (9 downto 0);
		y				: in signed (9 downto 0);
		
		cuadrante	: out unsigned (2 downto 0);
		radio			: out unsigned (9 downto 0)
		);
end component;

COMPONENT GENERADOR_PAREDES IS
	PORT(
		CLK		:	IN	STD_LOGIC;
		RAND		:	IN	STD_LOGIC_VECTOR(63 DOWNTO 0);
		MANTIENE	:	IN	STD_LOGIC;
		ADDR		:	IN	STD_LOGIC_VECTOR(5 DOWNTO 0);
		DATA		:	OUT	STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT PAREDES IS
	port(
		clk				:		in	std_logic;
		reset				:		in	std_logic;
		actualizar		:		in	std_logic;
		dificultad		:		in	std_logic_vector(1 downto 0);
		data				:		in	std_logic_vector(5 downto 0);
		cuadrante		:		in	unsigned(2 downto 0);
		radio				:		in	unsigned(9 downto 0);
		
		mantiene			:		out	std_logic;
		data_addr		:		out	std_logic_vector(5 downto 0);
		cuadrante_out	:		out	std_logic_vector(2 downto 0);
		visible			:		out	std_logic;
		isla				:		out	std_logic
	);
END COMPONENT;

component control_giro is 
port(
	clk					:	in	std_logic;
	reset					:	in	std_logic;
	Actualizar			:	in	std_logic;
	Random				:	in	std_logic_vector(63 downto 0);
	Subir_velocidad	:	in	std_logic;
	velocidad_prueba	:	out	unsigned(5 downto 0);
	angulo				:	out	unsigned(9 downto 0)
);
end component;

component Juego_Fsm is
	port(
		Clk				:	in	std_logic;
		Frame_inicio	:	in	std_logic;
		Frame_fin		:	in	std_logic;
		Nuevo_juego		:	in	std_logic;
		Colision			:	in	std_logic;
		Reset				:	in std_logic;
		
		Actualizar		:	out std_logic;
		Rst				:	out std_logic;
		Game_over		:	out std_logic	
	);
end component;

component CONTADOR is
	generic(max:integer:=16);
	port
	(
		-- Input ports
		Clk	: in  std_logic;
		EN		: in	std_logic;
		Rst	: in	std_logic;
		

		-- Output ports
		ovf: out std_logic
	);
end component;

component LFSR_64 is
	port
	(
		-- Input ports
		Clk	: in  std_logic;		
		Set	: in	std_logic;		
		En		: in	std_logic;

		-- Output ports
		b	: out std_logic_vector(63 downto 0)
	);
end component;

component senocoseno is
	port(
	clk		:	in	std_logic;
	angulo	:	in	unsigned(9 downto 0);
	seno		:	out	signed(11 downto 0);
	coseno	:	out	signed(11 downto 0)
	);
end component;

COMPONENT DIBUJO IS
	PORT(
		CLK		:	IN	STD_LOGIC;
		ALTERNA	:	IN	STD_LOGIC;
		CCOLOR	:	IN	STD_LOGIC;
		--RESET	:	IN	STD_LOGIC;
		DPAREDES	:	IN	STD_LOGIC;
		DISLA		:	IN	STD_LOGIC;
		DJUGADOR	:	IN	STD_LOGIC;
		CUADRANTE:	IN	STD_LOGIC_VECTOR(2 DOWNTO 0);
		RAND		:	IN	STD_LOGIC_VECTOR(63 DOWNTO 0);
		
		ROJO		:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		VERDE		:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		AZUL		:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
end component;

component jugador is
	port(
		Clk				: in	std_logic;
		Actualizar		: in	std_logic;
		Dificultad		: in	std_logic_vector(1 downto 0);
		Boton_der		: in	std_logic;
		Boton_izq		: in	std_logic;
		
		X_actual			: out	signed(9 downto 0);
		Y_actual			: out	signed(9 downto 0);
		X_anterior		: out	signed(9 downto 0);
		Y_anterior		: out	signed(9 downto 0)
	);
end component;

COMPONENT CIRCULO IS
	PORT(
		CLK	:	IN		STD_LOGIC;
		X1	:	IN		SIGNED(9 DOWNTO 0);	
		Y1	:	IN		SIGNED(9 DOWNTO 0);
		X2	:	IN		SIGNED(9 DOWNTO 0);
		Y2	:	IN		SIGNED(9 DOWNTO 0);
		
		DIBUJA:	OUT	STD_LOGIC
	);
END COMPONENT;

component Dificultad is
	port(
		Clk			:	in std_logic;
		switches		:	in	std_logic_vector(1 downto 0);
		gameover		:	in	std_logic;
		
		Dificultad	:	out std_logic_vector(1 downto 0);
		Leds_Rojo	:	out std_logic_vector(7 downto 0);
		Leds_Verde	:	out std_logic_vector(7 downto 0)
	);
end component;

component Compara_coordenadas is
	port(
		--inputs
		Xin1			: in signed(9 downto 0);
		Yin1			: in signed(9 downto 0);
		Xin2			: in signed(9 downto 0);
		Yin2			: in signed(9 downto 0);
	
		--outputs
		Comparacion		: out std_logic
	);
end component;

component FF_AND is
	port(
		Clk	: in	std_logic;
		IN1	: in	std_logic;
		IN2	: in	std_logic;
		
		OUT1	: out	std_logic
	);
end component;

COMPONENT PUNTAJE IS
	PORT(
		CLK			:	IN	STD_LOGIC;
		ACTUALIZAR	:	IN	STD_LOGIC;
		GAME_OVER	:	IN	STD_LOGIC;
		RESET			:	IN	STD_LOGIC;
		
		SEGUNDOS		:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
		SEGUNDOSX10	:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
		SEGUNDOSX100:	OUT	STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;
--------------------------------------------------------------------------------------------------------------------
END PACKAGE;
--------------------------------------------------------------------------------------------------------------------

PACKAGE BODY HexaPackage IS

function bit2bool(b: std_logic) return boolean is
begin
	if (b='1') then
		return true;
	else
		return false;
	end if;
end function bit2bool;

END PACKAGE BODY;