library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY SHIFT_REGISTER_RX IS
GENERIC(
	data_width:	integer:=8
	);
PORT(
	CLK:				IN		STD_LOGIC;
	RST:				IN		STD_LOGIC;
	DATAIN:			IN		STD_LOGIC;
	SHIFT:			IN		STD_LOGIC;
	DATAOUT:			OUT	STD_LOGIC_VECTOR(data_width-1 DOWNTO 0)
);
END SHIFT_REGISTER_RX;

ARCHITECTURE BEH OF SHIFT_REGISTER_RX IS
SIGNAL DATA:	STD_LOGIC_VECTOR(data_width-1 DOWNTO 0);
BEGIN
DATAOUT<=DATA;

SR: PROCESS (CLK, RST, SHIFT)
BEGIN
	IF(RST='1') THEN
		DATA<=(OTHERS=>'0');
	ELSIF(RISING_EDGE(CLK)) THEN
		IF (SHIFT='1') THEN
				DATA	<=	STD_LOGIC_VECTOR(UNSIGNED(DATA) SRL 1);
				DATA(data_width-1)	<= DATAIN;
		END IF;
	END IF;
END PROCESS;
END BEH;