library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY RS232_RX_FSM IS
	PORT(
		CLK:				IN	STD_LOGIC;
		RST:				IN	STD_LOGIC;
		TX:				IN	STD_LOGIC;
		
		SHIFT:			OUT	STD_LOGIC;
		DATA_OK:			OUT	STD_LOGIC
		);
END RS232_RX_FSM;

ARCHITECTURE BEH OF RS232_RX_FSM IS

SIGNAL CONT:		UNSIGNED(2 DOWNTO 0);
SIGNAL CONTCTRL:	STD_LOGIC_VECTOR(1 DOWNTO 0);	--00: NADA, 01: SUMA, 1X: RESETEA
TYPE STATE IS (IDLE, START, DATA, PARITY, STOP);
SIGNAL CS, NS: STATE;
BEGIN

NEXT_STATE:	PROCESS (CS, TX, CONT)
BEGIN
	CASE CS IS
		WHEN IDLE =>
			IF (TX='0') THEN
				NS <= DATA;
			ELSE
				NS <= IDLE;
			END IF;
		WHEN START => NS <= DATA;
		WHEN DATA =>
			IF (CONT = "111") THEN
				NS <= STOP;
			ELSE
				NS <= DATA;
			END IF;
		WHEN PARITY => NS <= STOP;
		WHEN STOP =>
			IF(TX='1') THEN
				NS <= IDLE;
			ELSE
				NS <= STOP;
			END IF;
		WHEN OTHERS => NS <= IDLE;
	END CASE;
END PROCESS;

CURRENT_STATE: PROCESS (CLK, RST)
BEGIN
	IF(RST='1') THEN
		CS <= IDLE;
	ELSIF(RISING_EDGE(CLK)) THEN
		CS <= NS;
	END IF;
END PROCESS;

OUTPUTS:	PROCESS (CS,RST,TX)
BEGIN
	IF (RST='1') THEN
		SHIFT	<='0';
		DATA_OK	<='0';
		CONTCTRL<="11";
	ELSE
		SHIFT	<='0';
		DATA_OK	<='0';
		CONTCTRL<="00";
		CASE CS IS
			WHEN IDLE => CONTCTRL<="11";
			WHEN START => NULL;
			WHEN DATA => 
				CONTCTRL<="01";
				SHIFT	<=	'1';
			--WHEN PARITY =>
				--SHIFT	<= '1';
			WHEN STOP =>
				IF(TX='1') THEN
					DATA_OK<='1';
				END IF;
			WHEN OTHERS => CONTCTRL<="11"; 
		END CASE;
	END IF;
END PROCESS;

COUNT_UP:	PROCESS (CLK,CONTCTRL)
BEGIN
	IF(RISING_EDGE(CLK)) THEN
		IF(CONTCTRL="01") THEN
			CONT<=CONT+1;
		ELSIF(CONTCTRL(1)='1') THEN
			CONT<="000";
		END IF;
	END IF;
END PROCESS;
END BEH;