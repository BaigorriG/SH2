library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
ENTITY CIRCULO IS
	PORT(
		CLK	:	IN		STD_LOGIC;
		X1	:	IN		SIGNED(9 DOWNTO 0);	
		Y1	:	IN		SIGNED(9 DOWNTO 0);
		X2	:	IN		SIGNED(9 DOWNTO 0);
		Y2	:	IN		SIGNED(9 DOWNTO 0);
		
		DIBUJA:	OUT	STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEH OF CIRCULO IS

CONSTANT	RADIO			:	SIGNED(9 DOWNTO 0)	:=	TO_SIGNED(2,10);
SIGNAL	DX,DY			:	SIGNED(9 DOWNTO 0);
BEGIN

CALCULA:PROCESS(CLK,DX,DY)
BEGIN
	IF RISING_EDGE(CLK) THEN
		DX<=X1-X2;		
		DY<=Y1-Y2;
		IF (DX*DX+DY*DY<RADIO*RADIO) THEN
			DIBUJA <= '1';
		ELSE 
			DIBUJA <= '0';
		END IF;
	END IF;
END PROCESS;

END ARCHITECTURE;